** sch_path: /foss/designs/prj_ADS1115_ic-1/design/design_comp/tb_comp_test.sch
**.subckt tb_comp_test
x1 VDD clk outn outp vin_p vin_n GND comp_test
V1 vin_p vin_n {vdiff}
V2 vin_n GND {vdd/2}
V3 clk GND dc 0 pulse(0, {vdd}, 1n, 50p, 50p, {per/2-1n}, {per})
V4 VDD GND {vdd}
**** begin user architecture code
 .lib cornerMOSlv.lib mos_tt


.param temp=27 vdd=1.5 per=1u vdiff=1m
.param Wnmos=1u Wpmos=2u
.param Lnmos=.3u Lpmos=.3u Lnmos2=1u
.option method=gear reltol=1e-5

.control
save all
tran 10p 4n
write tb_comp_test1.raw

alterparam vdiff=1u
;alterparam Wnmos=1u Wpmos=2u

reset
tran 10p 4n
write tb_comp_test2.raw
plot clk tran1.outp tran1.outn tran2.outp tran2.outn
.endc

**** end user architecture code
**.ends

* expanding   symbol:  comp_test.sym # of pins=7
** sym_path: /foss/designs/prj_ADS1115_ic-1/design/design_comp/comp_test.sym
** sch_path: /foss/designs/prj_ADS1115_ic-1/design/design_comp/comp_test.sch
.subckt comp_test VDD clk outn outp vin_p vin_n VSS
*.ipin clk
*.iopin VSS
*.iopin VDD
*.ipin vin_n
*.ipin vin_p
*.opin outn
*.opin outp
XM5p outn clk VDD VDD sg13_lv_pmos w=Wpmos l=Lpmos ng=1 m=1
XM4n outp outn VDD VDD sg13_lv_pmos w=Wpmos l=Lpmos ng=1 m=1
XM4p outn outp VDD VDD sg13_lv_pmos w=Wpmos l=Lpmos ng=1 m=1
XM5n outp clk VDD VDD sg13_lv_pmos w=Wpmos l=Lpmos ng=1 m=1
XM3p outn outp d2p VSS sg13_lv_nmos w=Wnmos l=Lnmos ng=1 m=1
XM3n outp outn d2m VSS sg13_lv_nmos w=Wnmos l=Lnmos ng=1 m=1
XM2n d2m clk d1m VSS sg13_lv_nmos w=Wnmos l=Lnmos ng=1 m=1
XM2p d2p clk d1p VSS sg13_lv_nmos w=Wnmos l=Lnmos ng=1 m=1
XM1n d1m vin_n VSS VSS sg13_lv_nmos w=Wnmos l=Lnmos2 ng=1 m=1
XM1p d1p vin_p VSS VSS sg13_lv_nmos w=Wnmos l=Lnmos2 ng=1 m=1
.ends

.GLOBAL GND
.end
