** sch_path: /foss/designs/prj_ADS1115_ic-1/design/design_comp/comp_test.sch
**.subckt comp_test out1m vdda pc out1p vinp vinm vssa
*.ipin clk
*.iopin vssa
*.iopin vdda
*.ipin vin_n
*.ipin vin_p
*.opin out1m
*.opin out1p
XM5p out1m clk vdda vdda sg13_lv_pmos w=Wpmos l=Lpmos ng=1 m=1
XM4n out1p out1m vdda vdda sg13_lv_pmos w=Wpmos l=Lpmos ng=1 m=1
XM4p out1m out1p vdda vdda sg13_lv_pmos w=Wpmos l=Lpmos ng=1 m=1
XM5n out1p clk vdda vdda sg13_lv_pmos w=Wpmos l=Lpmos ng=1 m=1
XM3p d2p out1p out1m vssa sg13_lv_nmos w=Wnmos l=Lnmos ng=1 m=1
XM3n d2m out1m out1p vssa sg13_lv_nmos w=Wnmos l=Lnmos ng=1 m=1
XM2n d1m clk d2m vssa sg13_lv_nmos w=Wnmos l=Lnmos ng=1 m=1
XM2p d1p clk d2p vssa sg13_lv_nmos w=Wnmos l=Lnmos ng=1 m=1
XM1n vssa vin_n d1m vssa sg13_lv_nmos w=Wnmos l=Lnmos ng=1 m=1
XM1p vssa vin_p d1p vssa sg13_lv_nmos w=Wnmos l=Lnmos ng=1 m=1
**.ends
.end
