** sch_path: /foss/designs/prj_ADS1115_ic-1/design/trail2-ota5.sch
**.subckt trail2-ota5 vdd vout ibias vinm vinp vss
*.ipin vss
*.ipin vdd
*.ipin ibias
*.ipin vinm
*.ipin vinp
*.opin vout
XM1 vout net1 vdd vdd sg13_lv_pmos w=0.22u l=0.3u ng=1 m=1
XM2 net2 vinm vout vss sg13_lv_nmos w=0.45u l=0.3u ng=1 m=1
XM3 net1 net1 vdd vdd sg13_lv_pmos w=0.22u l=0.3u ng=1 m=1
XM4 net2 vinp net1 vss sg13_lv_nmos w=0.45u l=0.3u ng=1 m=1
XM5 vss net3 net2 vss sg13_lv_nmos w=0.9u l=0.3u ng=1 m=1
XM6 vss net3 net4 vss sg13_lv_nmos w=0.9u l=0.3u ng=1 m=1
XM7 vss net3 net3 vss sg13_lv_nmos w=0.9u l=0.3u ng=1 m=1
XM8 net3 ibias ibias vdd sg13_lv_pmos w=0.44u l=0.3u ng=1 m=1
XM9 net4 ibias vdd vdd sg13_lv_pmos w=0.44u l=0.3u ng=1 m=1
**.ends
.end
